
module Lab2_sys (
	clk_clk,
	pio_data_seg_export,
	reset_reset_n);	

	input		clk_clk;
	output	[3:0]	pio_data_seg_export;
	input		reset_reset_n;
endmodule
